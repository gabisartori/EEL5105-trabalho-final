library ieee;
use ieee.std_logic_1164.all;

entity usertop is
port(

);
end usertop;

architecture rtl of usertop is
begin

end rtl;